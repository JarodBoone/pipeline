module opDecoder(control,regWrite,ALUOp,ALUSrc,memReg,branch,memWrite);
	input wire control; 
	
	// make these wires probably 
	output reg regWrite; 
	output reg ALUOp; 
	output reg ALUSrc; 
	output reg memReg; 
	output reg memWrite; 
	output reg branch; 


endmodule